module InstructionMemory(address, instruction, startin);

	input		  [31:0] address;
	input             startin;
	output reg [31:0] instruction;
	

	reg [7:0] m [67:0];

	always @(*) begin
	
		if(startin) begin
	/*		{m[0],m[1],m[2],m[3]} <= 32'b00100000000100000000000000000000;
			{m[4],m[5],m[6],m[7]} <= 32'b00100000000100010000000000000000;
			{m[8],m[9],m[10],m[11]} <= 32'b00100000000010000000000000101000;
			{m[12],m[13],m[14],m[15]} <= 32'b00010010000010000000000000000100;
			{m[16],m[17],m[18],m[19]} <= 32'b10001110000010010000000000000000;
			{m[20],m[21],m[22],m[23]} <= 32'b00000010001010011000100000100000;
			{m[24],m[25],m[26],m[27]} <= 32'b00100010000100000000000000000100;
			{m[28],m[29],m[30],m[31]} <= 32'b00001000000000000000000000000011;
			{m[32],m[33],m[34],m[35]} <= 32'b10101101000100010000000000000000;
			{m[36],m[37],m[38],m[39]} <= 32'b10001101000100100000000000000000;
			{m[40],m[41],m[42],m[43]} <= 32'b00001000000000000000000000001010;
			*/

			{m[0],m[1],m[2],m[3]} <=     32'b10001100000100000000000000000000; //Lw $s0, 0($0)
			{m[4],m[5],m[6],m[7]} <=     32'b10001100000100010000000000000100; //lw $s1, 4($0)
			{m[8],m[9],m[10],m[11]} <=   32'b10001100000100100000000000001000; //lw $s2, 8($0)
			{m[12],m[13],m[14],m[15]} <= 32'b10001100000100110000000000001100; //lw $s3, 12($0)
			{m[16],m[17],m[18],m[19]} <= 32'b00000000000000000000000000100000; // ADD $0, $0, $0
			{m[20],m[21],m[22],m[23]} <= 32'b00000000000000000000000000100000; // ADD $0, $0, $0
			{m[24],m[25],m[26],m[27]} <= 32'b00000000000000000000000000100000; // ADD $0, $0, $0
			{m[28],m[29],m[30],m[31]} <= 32'b00000000000000000000000000100000; // ADD $0, $0, $0
			{m[32],m[33],m[34],m[35]} <= 32'b00000010000100010100000000100000; //add $t0, $s0, $s1
			{m[36],m[37],m[38],m[39]} <= 32'b00000010010100110100100000100000; //add $t1, $s2, $s3
			{m[40],m[41],m[42],m[43]} <= 32'b00000001001010000101100000100000; //add $t3, $t1, $t0
			{m[44],m[45],m[46],m[47]} <= 32'b10101110000010110000000000101000; //sw $t3, 40($0)

		/*	{m[0],m[1],m[2],m[3]} <=     32'b00100000000010010000000000001010; 
			{m[4],m[5],m[6],m[7]} <=     32'b00000000000000000101000000100000; 
			{m[8],m[9],m[10],m[11]} <=   32'b00100000000010110000000000000001; 
			{m[12],m[13],m[14],m[15]} <= 32'b00000000000000000110000000100000; 
			{m[16],m[17],m[18],m[19]} <= 32'b00000000000000000111000000100000;
			{m[20],m[21],m[22],m[23]} <= 32'b00100000000011110000000000000100; 
			{m[24],m[25],m[26],m[27]} <= 32'b00010001001010100000000000001000; 
			{m[28],m[29],m[30],m[31]} <= 32'b00000001010010110101000000100000;  
			{m[32],m[33],m[34],m[35]} <= 32'b00000000000000000000000000100000; 
			{m[36],m[37],m[38],m[39]} <= 32'b10001101100011010000000000000000; 
			{m[40],m[41],m[42],m[43]} <= 32'b00000001110011010111000000100000; 
			{m[44],m[45],m[46],m[47]} <= 32'b00000001110010111000000000100000; 
			{m[48],m[49],m[50],m[51]} <= 32'b00000001110010111000100000100000; 
			{m[52],m[53],m[54],m[55]} <= 32'b00010000000000001111111111111000; 
			{m[56],m[57],m[58],m[59]} <= 32'b00000001100011110110000000100000; 
			{m[60],m[61],m[62],m[63]} <= 32'b00000000000000000000000000100000; 
			{m[64],m[65],m[66],m[67]} <= 32'b10101101100011100000000000000000; */

		end else begin
			
			instruction <= {m[address], m[address+1], m[address+2], m[address+3]};
		end
		
		
	end
		
endmodule


